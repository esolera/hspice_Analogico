** Profile: "_Fig1_12_MSD-_Fig1_12_MSD"  [ C:\Users\jbaker\Desktop\Ch1_MSD_PSpice\_Fig1_12_MSD\_fig1_12_msd-pspicefiles\_fig1_12_msd\_fig1_12_msd.sim ] 

** Creating circuit file "_Fig1_12_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC LIN 1000 10k 500Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig1_12_MSD.net" 


.END
