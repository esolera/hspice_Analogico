*** Figure 30.52 CMOS: Circuit Design, Layout, and Simulation ***

.tran 2n 2u 0 2n UIC

*#destroy all
*#run
*#let Vin=Vinsp-Vinsm
*#plot Vin
*#let Vout=Voutp-Voutm
*#plot Vout
*#plot Vout vs Vin 

*Input power and references
VDD VDD 0 DC 1
Vtrip Vtrip 0 DC 0.5
VCM VCM 0 DC 0.5
Vcip Vcip 0 DC 0 pwl 0 0 0.5u 0   0.501u 0.5 1.5u 0.5 1.501u 1
Vcim Vcim 0 DC 0 pwl 0 1 0.5u 1   0.501u 0.5 1.5u 0.5 1.501u 0

*Input Signal
Vinsp    Vinsp   0 DC 0 pulse 0.25 0.75 0 2u
Vinsm    Vinsm   0 DC 0 pulse 0.75 0.25 0 2u 

*Clock Signals
Vphi1  phi1  0 DC 0  Pulse 0 1   0    200p  200p  4n 10n
Vphi2  phi2  0 DC 0  Pulse 0 1   0    200p  200p  4n 10n
Vphi3  phi3  0 DC 0  Pulse 0 1   5n   200p  200p  4n 10n
R1 phi1 0 1MEG
R2 phi2 0 1MEG
R3 phi3 0 1MEG

*Use a VCVS for the op-amp
E1 Vopp VCM Vinp Vinm 100MEG
E2 VCM Vopm Vinp Vinm 100MEG

*Setup switched capacitors 
Cip Vinm Vbotip 1p 
Cfp Vinm Vbotfp 1p
Cim Vinp Vbotim 1p 
Cfm Vinp Vbotfm 1p

*Setup switches 
S1 Vbotfp Vinsp phi2 VTRIP switmod
S2 Vbotip Vinsp phi2 VTRIP switmod
S3 Vbotip Vcip   phi3 VTRIP switmod
S4 Vbotim Vcim   phi3 VTRIP switmod
S5 Vbotim Vinsm phi2 VTRIP switmod
S6 Vbotfm Vinsm phi2 VTRIP switmod
S7 Vopp Vbotfp  phi3 VTRIP switmod
S8 Vopp Vinm    phi1 VTRIP switmod
S9 Vopm Vinp    phi1 Vtrip switmod
S10 Vopm Vbotfm phi3 Vtrip switmod
S11 Vopp Voutp phi3 Vtrip  switmod
S12 Vopm Voutm phi3 Vtrip  switmod

Clp Voutp 0 10p
Clm Voutm 0 10p

.model switmod SW RON=1

.end
