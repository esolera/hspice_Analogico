** Profile: "SCHEMATIC1-_Fig2_40_mismatch_MSD"  [ c:\users\homepc\documents\spring 2013\pspice_cmosedu\msd\ch2_msd_pspice\_fig2_40_mismatch_msd\_fig2_40_mismatch_msd-pspicefiles\schematic1\_fig2_40_mismatch_msd.sim ] 

** Creating circuit file "_Fig2_40_mismatch_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500ns 0 .01n SKIPBP 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
