*** Figure 1.21 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vin vout

.tran 10u 16m 

Vin	Vin	0	DC	0	SIN 0 1 200
R1	Vin	Vout	1k
CL	Vout	0	1u

.end
