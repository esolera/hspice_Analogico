*** Figure 2.23 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vin vout

.tran 100p 100n 

O1	Vin	0	Vout	0	TRC
Rload	Vout	0	1G
Vin	vin	0	DC	0	pulse 0 1 5n 0

.model TRC 	ltra	R=5k 	C=5f	len=50

.end
