** Profile: "Fig2_19-diode"  [ C:\Users\jbaker\Desktop\PSpice_CMOSedu\Chap2_PSpice\Fig2_19\Fig2_19-pspicefiles\Fig2_19\diode.sim ] 

** Creating circuit file "diode.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig2_19-pspicefiles/Fig2_19.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 25ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig2_19.net" 


.END
