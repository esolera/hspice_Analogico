** Profile: "_Fig3_48_MSD-_Fig3_48_MSD"  [ C:\Users\jbaker\Desktop\Ch3_MSD_PSpice\_fig3_48_msd-pspicefiles\_fig3_48_msd\_fig3_48_msd.sim ] 

** Creating circuit file "_Fig3_48_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5us 0 .01u SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig3_48_MSD.net" 


.END
