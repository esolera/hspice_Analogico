*** Figure 30.36 CMOS: Circuit Design, Layout, and Simulation ***

.tran 2n 500n 0 2n UIC

*#destroy all
*#run
*#plot Vopp Vopm Vinsp
*#plot Vinm Vinp

*Input power and references
VDD VDD 0 DC 1
Vtrip Vtrip 0 DC 0.5
VCM VCM 0 DC 0.5

*Input Signal
Vinsp    Vinsp   0 DC 0 Sin 0.5 0.5 2.5MEG
Vinsm    Vinsm   0 DC 0.5

*Clock Signals
Vphi1  phi1  0 DC 0  Pulse 0 1   0    200p  200p  4n 10n
Vphi2  phi2  0 DC 0  Pulse 0 1   0    200p  200p  4n 10n
Vphi3  phi3  0 DC 0  Pulse 0 1   5n   200p  200p  4n 10n
R1 phi1 0 1MEG
R2 phi2 0 1MEG
R3 phi3 0 1MEG

*Use a VCVS for the op-amp
E1 Vopp VCM Vinp Vinm 100MEG
E2 VCM Vopm Vinp Vinm 100MEG

*Setup switched capacitors  
Cfp Vinm Vbotfp 0.9p 
Cfm Vinp Vbotfm 1p

*Setup switches 
S1 Vbotfp Vinsp phi2 VTRIP switmod
S6 Vbotfm Vinsm phi2 VTRIP switmod
S7 Vopp Vbotfp  phi3 VTRIP switmod
S8 Vopp Vinm    phi1 VTRIP switmod
S9 Vopm Vinp    phi1 Vtrip switmod
S10 Vopm Vbotfm phi3 Vtrip switmod

.model switmod SW RON=1

.end
