*** Figure 23.14 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#set temp=0
*#run
*#set temp=25
*#run
*#set temp=50
*#run
*#set temp=75
*#run
*#set temp=100
*#run
*#plot dc1.i(vdd) dc2.i(vdd) dc3.i(vdd) dc4.i(vdd) dc5.i(vdd)
*#plot dc1.vref dc2.vref dc3.vref dc4.vref dc5.vref

.option scale=50n
.dc VDD 0 1.2 1m

VDD 	VDD	0	DC	1 

M1	Vbiasn	Vbiasn	0	0	N_50n L=2 W=10
M2	Vref	Vref	Vr	0	N_50n L=2 W=40
M3	Vbiasn	Vbiasp	VDD	VDD	P_50n L=2 W=100
M4	Vref	Vbiasp	VDD	VDD	P_50n L=2 W=100

Rbias	Vr	0	5.5k 	Rmod
.model RMOD R TC1=0.002

*amplifier 
MA1	Vamp	Vref	0	0	N_50n L=2 W=10
MA2	Vbiasp	Vbiasn	0	0	N_50n L=2 W=10
MA3	Vamp	Vamp	VDD	VDD	P_50n L=2 W=100
MA4	Vbiasp	Vamp	VDD	VDD	P_50n L=2 W=100

*start-up stuff
MSU1	Vsur	Vbiasn	0	0	N_50n L=2   W=10
MSU2	Vsur	Vsur	VDD	VDD	P_50n L=20  W=10
MSU3	Vbiasp	Vsur	Vbiasn	0	N_50n L=1   W=10

.include cmosedu_models.txt  

.end
   

