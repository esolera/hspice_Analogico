** Profile: "fig2-23-diode"  [ C:\USERS\student\Desktop\Chap2_PSpice\Fig2-23\Fig2_23-PSpiceFiles\fig2-23\diode.sim ] 

** Creating circuit file "diode.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../fig2_23-pspicefiles/fig2_23.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\fig2-23.net" 


.END
