** Profile: "Tab9_1_ftp-ac"  [ C:\Users\jbaker\Desktop\Chap9_PSpice\Tab9_1_ftp\Tab9_1_ftp-pspicefiles\Tab9_1_ftp\ac.sim ] 

** Creating circuit file "ac.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Tab9_1_ftp-pspicefiles/Tab9_1_ftp.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10MEG 10G
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Tab9_1_ftp.net" 


.END
