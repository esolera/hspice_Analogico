*** Figure 30.9 CMOS: Circuit Design, Layout, and Simulation ***

.tran 1n 640n 10n 1n UIC

*#destroy all
*#run
*#let bin5=b5+7.5
*#let bin4=b4+6
*#let bin3=b3+4.5
*#let bin2=b2+3
*#let bin1=b1+1.5 
*#let bin0=b0+0
*#plot bin5 bin4 bin3 bin2 bin1 bin0
*#plot out ylimit .48 .52 xlimit 10n 600n

VDD VDD 0 DC 1
VREFP VREFP 0 DC 1
VREFM VREFM 0 DC 0.0

VB5 B5 0 DC 0 pulse 1 0 0 200p 200p 319.8n  640n
VB4 B4 0 DC 0 pulse 1 0 0 200p 200p 159.8n  320n
VB3 B3 0 DC 0 pulse 1 0 0 200p 200p 79.8n   160n
VB2 B2 0 DC 0 pulse 1 0 0 200p 200p 39.8n   80n
VB1 B1 0 DC 0 pulse 1 0 0 200p 200p 19.8n   40n
VB0 B0 0 DC 0 pulse 1 0 0 200p 200p 9.8n    20n

*Generate Logic switching point, or trip, voltage
R1 VDD trip 100MEG
R2 trip 0   100MEG

*Make resistive ladder
R11 Vrefp out 10k
R12 Vrefm out 10k
R22 out outl 100k
X5 trip B5 in5 outl Vrefp Vrefm R2R
X4 trip B4 in4 in5 Vrefp Vrefm R2R
X3 trip B3 in3 in4 Vrefp Vrefm R2R
X2 trip B2 in2 in3 Vrefp Vrefm R2R
X1 trip B1 in1 in2 Vrefp Vrefm R2R
X0 trip B0 in0 in1 Vrefp Vrefm R2R
RT in0 0 10k

.subckt R2R trip BX in out Vrefp Vrefm
SH 	Vrefp	2R	BX	trip 	Switmod
SL	Vrefm	2R	trip	BX	Switmod
R2R	2R	out	20k
R1R	out	in	10k	
.model switmod SW
.ends

.end
