*** Figure 23.5 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#set temp=0
*#run
*#set temp=25
*#run
*#set temp=50
*#run
*#set temp=75
*#run
*#set temp=100
*#run
*#plot dc1.vref dc2.vref dc3.vref dc4.vref dc5.vref

.option scale=1u
.dc VDD 4 6 1m

VDD 	VDD	0	DC	5
R1	VDD	VREF	10k	RMOD
M1	VREF	VREF	0	0	N_1u L=2 W=10

.model RMOD R TC1=0.002

.include cmosedu_models.txt

.end
      