*** Example 8.10 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot onoise_spectrum 
*#print all

.noise	 V(Vout,0)	Vs 	dec  	100 	1 	1k 
Rs	 Vs 	Vout 	10k 
Gin	 Vout 	0 	Vout 	0 	1e-3 
Vs	 Vs 	0	dc 	0 	ac 	1
.print noise all
.end