*** Figure 1.31 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vout

.tran 100p 8n UIC

Vclk	clk	0	pulse -1 1 2n

Vin	Vin	0	DC	5
R1	Vin	Vouts	1k
S1	Vouts	Vout	0	clk	switmodel
R2	Vout	0	1k
L1	Vout	0	10u 	IC=5mA

.model switmodel sw ron=0.1 

.end
