*** Figure 1.10 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#print all

.op

Vin	1	0	DC	1
R1	1	2	1k
R2	2	0	2k

.end