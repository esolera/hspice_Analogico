** Profile: "_Fig3_28_MSD_alt-_Fig3_28_MSD_alt"  [ C:\Users\jbaker\Desktop\Ch3_MSD_PSpice\_fig3_28_msd_alt-pspicefiles\_fig3_28_msd_alt\_fig3_28_msd_alt.sim ] 

** Creating circuit file "_Fig3_28_MSD_alt.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 10k 200meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig3_28_MSD_alt.net" 


.END
