*** SPICE Circuit File of 3TO1_DIV_LAY  02/27/04 09:58:43

* Start of C:\Lasi7\Mosis\3to1_div.txt

*#destroy all
*#run
*#plot vin vout

.dc vin 0 1 1m

vin vin 0 DC 0
* End of C:\Lasi7\Mosis\3to1_div.txt

* MAIN 3TO1_DIV_LAY
R1 Vin Vout 2k
R2 vn1 Vout 2k
R3 vn1 0 2k
.END
