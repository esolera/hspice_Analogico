*** Figure 4.6 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vin vout1 
*#plot vin vout2 xlimit 40p 140p

.tran 1p 2500p 

Vin	vin	0	DC	0	pulse 0 1 50p 0

O1	Vin	0	Vout1	0	poly_nosilicide
Rload1	Vout1	0	1G

O2	Vin	0	Vout2	0	poly_silicide
Rload2	Vout2	0	1G

.model 	poly_nosilicide ltra	R=200 	C=9e-18 len=1000

.model 	poly_silicide 	ltra	R=5 	C=9e-18 len=1000
.end
