*** Figure 14.2 (PMOS) CMOS: Circuit Design, Layout, and Simulation *** 

*#destroy all
*#run
*#let ID=-i(vdd)
*#plot log(ID)

.option scale=50n
.dc	vsg	-0.1	1	1m

vdd	vdd	0	DC	1
vsg	vdd	vsg	DC	0

M1	0	vsg	vdd	vdd	P_50n L=1 W=10

.include cmosedu_models.txt 

.end
   

