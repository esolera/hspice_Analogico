*** Figure 20.26 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#set temp=0
*#run
*#set temp=27
*#run
*#set temp=100
*#run
*#let Iref0=-tran1.VDD#branch
*#let Iref27=-tran2.VDD#branch
*#let Iref100=-tran3.VDD#branch
*#plot Iref0 Iref27 Iref100

.option scale=50n
.tran 1m 1

VDD	VDD	0 	DC 	1

R1	VD1	0	65k	RMOD
M1	VD1	VD1	VDD	VDD	P_50n L=2 W=100

.model RMOD R TC1=0.002

.include cmosedu_models.txt

.end
   

