** Profile: "SCHEMATIC1-_Fig1_25_K_is_4_AC_MSD"  [ C:\Users\HomePC\Documents\Spring 2013\CMOSEDU_PSPICE\MSD\Ch1_MSD_Pspice\_Fig1_25_K_is_4_AC_MSD-PSpiceFiles\SCHEMATIC1\_Fig1_25_K_is_4_AC_MSD.sim ] 

** Creating circuit file "_Fig1_25_K_is_4_AC_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC LIN 1000 1k 100MEG
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
