*** Figure 9.30 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#set temp=0
*#run
*#set temp=50
*#run
*#set temp=100
*#run
*#plot -dc1.vds#branch -dc2.vds#branch -dc3.vds#branch ylimit 10u 50u xlimit 0.25 0.45
*#plot -dc1.vds#branch -dc2.vds#branch -dc3.vds#branch ylimit 0 600u


.option scale=50n
.DC 	VGS	0	1	1m

VDS 	VDS	0	DC	1
VGS	VGS	0	DC	0

M1	VDS	VGS	0	0	N_50n L=2 W=50

.include cmosedu_models.txt

.end
   
