** Profile: "_Fig2_48_MSD-_Fig2_48_MSD"  [ C:\Users\jbaker\Desktop\Ch2_MSD_Pspice\_Fig2_48_MSD\_Fig2_48_MSD-pspicefiles\_Fig2_48_MSD\_Fig2_48_MSD.sim ] 

** Creating circuit file "_Fig2_48_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500ns 0 .01n SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig2_48_MSD.net" 


.END
