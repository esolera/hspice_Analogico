*** Figure 9.29 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#set temp=0
*#run
*#set temp=50
*#run
*#set temp=100
*#run
*#plot -dc1.vds#branch -dc2.vds#branch -dc3.vds#branch 


.option scale=1u
.DC 	VGS	0.8	1.6	1m

VDS 	VDS	0	DC	2
VGS	VGS	0	DC	0

M1	VDS	VGS	0	0	N_1u L=2 W=10
                                                                     
.include cmosedu_models.txt

.end
      
