*** Figure 1.13 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#print all

.TF 	V(Vout,0) Vin

Vin	Vin	0	DC	1
R1	Vb	0	3k
R2	Vt	Vout	1k
R3	Vout	0	2k
E1	vt	vb	Vin	0	23

.end