*** Figure 9.24 (NMOS) CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#let ID=-VDD#branch
*#plot ID
*#let ro=1/deriv(ID)
*#plot ro

.option scale=1u
.dc VDD 0 5 1m

VDD 	VDD	0	DC	5
VGN	VGN	0	DC	1.05

MN	VDD	VGN	0	0	N_1u L=2 W=10

.include cmosedu_models.txt  

.end
      