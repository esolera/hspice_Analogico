*** Example 8.6 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot onoise_spectrum xlog
*#print all

.noise	 V(Vout,0) 	Vin 	dec  	100 	1 	1G 
R1	 Vin 		Vout 	10k 
C1	 Vout 	0 	1p 
Vin	 Vin 	0	dc 	0 	ac 	1
.print noise all	
.end