** Profile: "Fig9_34_PMOS-ac"  [ C:\Users\jbaker\Desktop\Chap9_PSpice\Fig9_34_PMOS\fig9_34_pmos-pspicefiles\fig9_34_pmos\ac.sim ] 

** Creating circuit file "ac.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../fig9_34_pmos-pspicefiles/fig9_34_pmos.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10meg 10G
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig9_34_PMOS.net" 


.END
