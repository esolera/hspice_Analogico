** Profile: "Fig5_2-dc"  [ C:\Users\jbaker\Desktop\PSpice_CMOSedu\Chap5_PSpice\Fig5_2\Fig5_2-pspicefiles\Fig5_2\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig5_2-pspicefiles/Fig5_2.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_Vr 0.9 1.1 0.01 
.TEMP 0 27 100
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig5_2.net" 


.END
