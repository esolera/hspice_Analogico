*** Figure 29.48 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vin vout_digital vout_filtered


Vin Vin 0 0.4
Vphi1 phi1 0 PULSE(0 5 0 200p 200p 4n 10n)
VDD VDD 0 5
CF N001 vointeg 1p
CI N003 N002 1p
Vphi2 phi2 0 PULSE(0 5 5n 200p 200p 4n 10n)
XX4 vointeg 0 N004 VDD phi1 ideal_clocked_comparator
XX1 N001 0 vointeg op_amp
XX2 N003 N001 phi2 VDD switch_1
XX3 Vin N002 phi1 VDD switch_1
XX7 N003 0 phi1 VDD switch_1
XX8 N002 Vout_digital phi2 VDD switch_1
XX5 VREFP Vout_digital N005 VDD switch_1
XX9 N004 N005 VDD inverter
XX10 Vout_digital VREFM N004 VDD switch_1
R1 Vout_digital Vout_filtered 10k
C1 Vout_filtered 0 10p
VREFP VREFP 0 1
VREFM VREFM 0 -1

* block symbol definitions
.subckt ideal_clocked_comparator Vinm Vinp Vout VDD Clock
S1 Vout VDD N001 0 switmod
S2 0 Vout 0 N001 switmod
XX1 N002 N001 Clock VDD sample_and_hold
E1 N002 0 Vinp Vinm 1
.model switmod SW
.ends ideal_clocked_comparator

.subckt op_amp Vinm Vinp Out
G1 0 Out Vinp Vinm 1000
R1 Out 0 1
.ends op_amp

.subckt switch_1 P1 P2 clk VDD
S1 P2 P1 clk Vtrip switmod
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
.model switmod SW
.ends switch_1

.subckt inverter In Out VDD
S3 Out VDD N001 In switmod
S4 0 Out In N001 switmod
E1 N001 0 VDD 0 0.5
.model switmod SW
.ends inverter

.subckt sample_and_hold Vin Outsh Clock VDD
S1 Vins Vinb Vtrip Clock switmod
C1 Vins 0 1e-10
S2 N001 Vins clock Vtrip switmod
C2 N001 0 1e-16
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
Ebufout Outsh 0 N001 0 1
Ebufin Vinb 0 Vin 0 1
.model switmod SW
.ends sample_and_hold

.tran 0 500n 0 2n uic
* Nonoverlapping clocks
.options plotwinsize=0

.end

