** Profile: "SCHEMATIC1-_Fig3_23_MSD"  [ C:\USERS\HOMEPC\DOCUMENTS\SPRING 2013\PSPICE_CMOSEDU\MSD\CH3_MSD_PSPICE\_FIg3_23_MSD-PSpiceFiles\SCHEMATIC1\_Fig3_23_MSD.sim ] 

** Creating circuit file "_Fig3_23_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2000ns 0 .01n SKIPBP 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
