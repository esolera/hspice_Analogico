*** Figure 11.11 with Varying load C from
*** CMOS: Circuit Design, Layout, and Simulation


*#destroy all
*#let cap = 25f
*#while cap <= 100f
*#    alter @Cload[capacitance] = cap
*#    run
*#    let cap = cap + 25f
*#end
** plot load C from 25f to 100f
*#plot tran1.vout tran2.vout tran3.vout tran4.vout vin

.option scale=50n
.tran 10p 2n UIC

vdd	vdd	0	DC	1
Vin	vin	0	DC	0	pulse 0 1 500p 0 0 1n 2n

M1	vout	vin	0	0	N_50n L=1 W=10	
M2	vout	vin	vdd	vdd	P_50n L=1 W=20

Cload	vout	0	50f	

.include cmosedu_models.txt 

.end
   

