*** Equation 21.75 NOISE CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run

* Plot PSD's of the amplifier's input and output noise 
*#plot inoise_spectrum loglog
*#plot onoise_spectrum loglog

* Print the RMS input and output noise voltages
*#let VonoiseRMS=sqrt(onoise_total)
*#let VinoiseRMS=sqrt(inoise_total)
*#print vonoiseRMS VinoiseRMS

.noise	 v(Vout,0)	Vin 	dec  	100 	1 	100MEG 
.options scale=50n

VDD	VDD	0	DC	1
Vin	Vin	0	DC	350m	AC	1

* Bias the MOSFETs at the operating points in Table 9.2 (back inside cover)

M2	Vout	VACGND	VDD	VDD	P_50n L=2 W=100
RBIG	VACGND	Vout	100MEG
CBIG	VACGND	0	1u
M1	Vout	Vin	0	0	N_50n L=2 W=50


.include cmosedu_models.txt  

.end
   

