*** Figure 9.27 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#let ID=-VDS#branch
*#let gm=deriv(ID)
*#plot gm
*#plot ID

.option scale=50n
.DC 	VGS	0	1	1m

VDS 	VDS	0	DC	.1
VGS	VGS	0	DC	0

M1	VDS	VGS	0	0	N_50n L=2 W=10

.include cmosedu_models.txt


.end
   
