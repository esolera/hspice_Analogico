*** Figure 30.58 CMOS: Circuit Design, Layout, and Simulation ***

.tran .2n 200n 50n .2n UIC

*#destroy all
*#run
*#plot phi1+2.5 phi2+1.25 phi3
*#let error=1-Voutp
*#plot error ylimit 0 10m

*Input power and references
VDD VDD 0 DC 1
Vtrip Vtrip 0 DC 0.5
VCM VCM 0 DC 0.5
Vcip Vcip 0 DC 0.5 
Vcim Vcim 0 DC 0.5 

*Input Signal
Vinsp    Vinsp   0 DC 1.0
Vinsm    Vinsm   0 DC 0.5

*Clock Signals
Vphi1  phi1  0 DC 0  Pulse 0 1   0    200p  200p  4n 10n
Vphi2  phi2  0 DC 0  Pulse 0 1   0    200p  200p  4n 10n
Vphi3  phi3  0 DC 0  Pulse 0 1   5n   200p  200p  4n 10n
R1 phi1 0 1MEG
R2 phi2 0 1MEG
R3 phi3 0 1MEG

*Use a VCVS for the op-amp
E1 Vopp VCM Vinp Vinm 100MEG
E2 VCM Vopm Vinp Vinm 100MEG

*Setup switched capacitors 
Cip Vinm Vbotip 1.00p 
Cfp Vinm Vbotfp 1.02p
Cim Vinp Vbotim 1.04p 
Cfm Vinp Vbotfm 1.06p

*Setup switches 
S1 Vbotfp Vinsp  phi2 VTRIP  switmod
S2 Vbotip Vinsp  phi2 VTRIP  switmod
S3 Vbotip Vcip   phi3 VTRIP  switmod
S4 Vbotim Vcim   phi3 VTRIP  switmod
S5 Vbotim Vinsm  phi2 VTRIP  switmod
S6 Vbotfm Vinsm  phi2 VTRIP  switmod
S7 Vopp Vbotfp   phi3 VTRIP  switmod
S8 Vopp Vinm     phi1 VTRIP  switmod
S9 Vopm Vinp     phi1 Vtrip  switmod
S10 Vopm Vbotfm  phi3 Vtrip  switmod
S11 Vopp Voutp   phi3 Vtrip  switmod
S12 Vopm Voutm   phi3 Vtrip  switmod

Clp Voutp 0 10p
Clm Voutm 0 10p

.model switmod SW RON=1

.end
