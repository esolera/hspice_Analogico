** Profile: "Fig10_5_NMOS-dc"  [ C:\Users\jbaker\Desktop\Chap10_PSpice\Fig10_5_NMOS\Fig10_5_nmos-pspicefiles\Fig10_5_nmos\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig10_5_nmos-pspicefiles/Fig10_5_nmos.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VDS 0 5 1m 
+ LIN V_VGS 0 5 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig10_5_NMOS.net" 


.END
