*** Figure 21.14 NOISE CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run

* Plot PSD's of the amplifier's input and output noise 
*#plot inoise_spectrum loglog
*#plot onoise_spectrum loglog

* Noting that the gain of this amplifier is around 1 so input and output noise are equal
*#print inoise_total onoise_total

* Print the RMS input and output noise voltages
*#let VonoiseRMS=sqrt(onoise_total)
*#let VinoiseRMS=sqrt(inoise_total)
*#print vonoiseRMS VinoiseRMS

.noise	 v(Vout,0)	Vin 	dec  	100 	1 	100MEG 
.options scale=50n

VDD	VDD	0	DC	1
Vin	Vin	0	DC	350m	AC	1

* Bias the MOSFETs at the operating points in Table 9.2 (back inside cover)

M2	Vout	Vout	VDD	VDD	P_50n L=2 W=100
M1	Vout	Vin	0	0	N_50n L=2 W=50


.include cmosedu_models.txt    

.end
   

