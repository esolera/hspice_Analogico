*** Figure 1.12 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#print all

.TF 	I(Vmeas) Vin

Vin	Vin	0	DC	1
R1	Vin	Vout	1k
R2	Vout	Vmeas	2k
Vmeas	Vmeas	0	DC	0

.end