*** Example 8.18 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot onoise_spectrum 
*#print all

.noise	V(Vout,0)	Vplus 	dec  	100 	1 	1000G 

Vplus	Vplus	0	dc	0	ac	1
Rf	Vout	Vminus	100k
Cf	Vout	Vminus 	1000pf
Eopamp	Vout	0	Vplus	Vminus 100MEG

.print noise all
.end