** Profile: "Ex8_5-noise"  [ C:\Users\jbaker\Desktop\PSpice_CMOSedu\Chap8_PSpice\Ex8_5\Ex8_5-pspicefiles\Ex8_5\noise.sim ] 

** Creating circuit file "noise.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100 1 1k
.NOISE V([VOUT],[0]) V_Vin 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Ex8_5.net" 


.END
