** Profile: "Fig9_24_NMOS-dc"  [ C:\Users\jbaker\Desktop\Chap9_PSpice\Fig9_24_NMOS\Fig9_24_nmos-pspicefiles\Fig9_24_nmos\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig9_24_nmos-pspicefiles/Fig9_24_nmos.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VDS 0 5 0.005 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig9_24_NMOS.net" 


.END
