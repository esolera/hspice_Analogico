*** Figure 9.8 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#let VGS4=VG3-VD2
*#plot VD2 VGS4

.option scale=1u
.dc 	Iinject	-1u 	1u 	10n	

VDD 	VDD	0	DC	5
Ibias	VDD	VG3	DC	1u
Iinject	0	VD2	DC	0

M1	VG1	VG1	0	0	N_1u L=1 W=10
M2	VD2	VG1	0	0	N_1u L=1 W=10
M3	VG3	VG3	VG1	0	N_1u L=1 W=10
M4	VDD	VG3	VD2	0	N_1u L=1 W=10

.inculde cmosedu_models.txt 

.end
      