*** Example 8.13 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot onoise_spectrum 
*#print all

.noise	V(Vout,0)	Vs 	dec  	100 	1 	1000G 

Vs	Vs	0	dc	1.7	ac	1
Rs	Vs	Vout	1k
D1	0 	Vout 	Diode

.model Diode D TT=10n Rs=0 cj0=25e-15 vj=1 m=.5
.print noise all
.end