*** Figure 14.2 CMOS: Circuit Design, Layout, and Simulation *** 

*#destroy all
*#run
*#let ID=-i(vdd)
*#plot log(ID)

.option scale=50n
.dc	vgs	-0.1	1	1m

vdd	vdd	0	DC	1
vgs	vgs	0	DC	0

M1	vdd	vgs	0	0	N_50n L=1 W=10

.include cmosedu_models.txt 

.end
   

