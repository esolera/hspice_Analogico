*** Figure 18.26 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot V1 V1out
*#plot V2 V2out

.option scale=50n
.tran	.1n 100n

V1	V1	0	DC	0	PULSE 0 1 0 0 0 4n 20n
R1	V1	V1out	1k
C1	V1out	0	10p


V2	V2	0	DC	0	PULSE 0 1 0 0 0 12n 20n
R2	V2	V2out	1k
C2	V2out	0	10p

.include cmosedu_models.txt 

.end
   
