*** Figure 28.21 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot Qe_no_error Qe_error

Vclock clk 0 PULSE(0 1 5n 100p 100p 4.9n 10n)
VDD VDD 0 1
Vin Vin 0 PULSE(0 1 0 10u)
XX2 b2 b1 b0 Vout_error VDD 0 VDD ideal_3_bit_dac
Eqe Qe_error 0 Vout_error Vin 1
XX1 b2 b1 b0 Vin VDD 0 clk VDD error_3_bit_adc
XX3 N001 N002 N003 Vout VDD 0 VDD ideal_3_bit_dac
Eqe1 Qe_no_error 0 Vout Vin 1
XX4 N001 N002 N003 Vin VDD 0 clk VDD ideal_3_bit_adc

* block symbol definitions
.subckt ideal_3_bit_dac B2 B1 B0 Vout Vrefp Vrefm VDD
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
S7 B2L Vone B2 Vtrip switmod
S8 0 B2L Vtrip B2 switmod
S13 B1L Vone B1 Vtrip switmod
S14 0 B1L Vtrip B1 switmod
S15 B0L Vone B0 Vtrip switmod
S16 0 B0L Vtrip B0 switmod
B1 Vout 0 V=((v(vrefp)-v(vrefm))/8)*(v(B2L)*4+v(B1L)*2+v(B0L))+v(vrefm)
R3 Vrefp Vrefm 100MEG
Vone Vone 0 1
.model switmod SW
.ends ideal_3_bit_dac

.subckt error_3_bit_adc B2 B1 B0 Vin Vrefp Vrefm Clock VDD
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
B1 VCM 0 V=(V(VREFP)-V(VREFM))/2
BPIP PIPIN 0 V=V(OUTSH)-V(VREFM)+((V(VREFP)-V(VREFM))/16)
XU8 VDD Vtrip VCM N001 B1 N002 adcbit
XU9 VDD Vtrip VCM N002 B0 NC_01 adcbit
XU10 Vin OUTSH clock VDD sample_and_hold
XX1 VDD Vtrip VCM PIPIN B2 N001 error_adcbit
.ends error_3_bit_adc

.subckt ideal_3_bit_adc B2 B1 B0 Vin Vrefp Vrefm Clock VDD
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
B1 VCM 0 V=(V(VREFP)-V(VREFM))/2
BPIP PIPIN 0 V=V(OUTSH)-V(VREFM)+((V(VREFP)-V(VREFM))/16)
XU7 VDD Vtrip VCM PIPIN B2 N001 adcbit
XU8 VDD Vtrip VCM N001 B1 N002 adcbit
XU9 VDD Vtrip VCM N002 B0 NC_01 adcbit
XU10 Vin OUTSH clock VDD sample_and_hold
.ends ideal_3_bit_adc

.subckt adcbit VDD Vtrip VCM Vin Bitout Vout
S3 Bitout VDD Vin VCM switmod
S4 0 Bitout VCM Vin switmod
S5 Vout Vinh Bitout Vtrip switmod
S6 Vinl Vout Vtrip Bitout switmod
E1 Vinh 0 Vin VCM 2
E2 Vinl 0 Vin 0 2
.model switmod SW
.ends adcbit

.subckt sample_and_hold Vin Outsh Clock VDD
S1 Vins Vinb Vtrip Clock switmod
C1 Vins 0 1e-10
S2 N001 Vins clock Vtrip switmod
C2 N001 0 1e-16
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
Ebufout Outsh 0 N001 0 1
Ebufin Vinb 0 Vin 0 1
.model switmod SW
.ends sample_and_hold

.subckt error_adcbit VDD Vtrip VCM Vin Bitout Vout
S3 Bitout VDD Vin VCM switmod
S4 0 Bitout VCM Vin switmod
S5 Vout Vinh Bitout Vtrip switmod
S6 Vinl Vout Vtrip Bitout switmod
E1 Vinh 0 Vin VCM 2.5
E2 Vinl 0 Vin 0 1.9
.model switmod SW
.ends error_adcbit

.tran 0 10u 0 .1n uic
.options plotwinsize=0

.end
