*** Figure 29.23_V2 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vout vin

*** CELL: Ideal_Differencer_1{sch}
.SUBCKT Ideal_Differencer_1 im ip om op

* Spice Code nodes in cell cell 'Ideal_Differencer_1{sch}'
E  op  om  ip  im  1
.ENDS Ideal_Differencer_1

*** CELL: Ideal_Switch{sch}
.SUBCKT Ideal_Switch contrlm contrlp in out

* Spice Code nodes in cell cell 'Ideal_Switch{sch}'
Sswitch  in out  contrlp contrlm  switmod
.model switmod sw
.ENDS Ideal_Switch

*** CELL: Ideal_Opamp{sch}
.SUBCKT Ideal_Opamp Vm Vo Vp
** GLOBAL gnd
Rres@0 Vp Vm 1410.065meg
Rres@1 Vo gnd 1

* Spice Code nodes in cell cell 'Ideal_Opamp{sch}'
G1 Vo 0  Vp  Vm 100MEG
.ENDS Ideal_Opamp

*** CELL: Ideal_Sample&Hold{sch}
.SUBCKT Ideal_Sample_Hold Vclk Vin Voutsh vdd
** GLOBAL gnd
Ccap@0 gnd Vins 0.1n
Ccap@1 gnd net@32 0.1f
Rres@0 vdd Vtrip 100000k
Rres@1 Vtrip gnd 100000k
XIdeal_sw@0 Vclk Vtrip Vinb Vins Ideal_Switch
XIdeal_sw@1 Vtrip Vclk Vins net@32 Ideal_Switch
Xideal_op@0 Voutsh Voutsh net@32 Ideal_Opamp
Xideal_op@1 Vinb Vinb Vin Ideal_Opamp
.ENDS Ideal_Sample_Hold

*** CELL: Ideal_clocked_comparator{sch}
.SUBCKT Ideal_clocked_comparator Clock Vinm Vinp Vout vdd
** GLOBAL gnd
XIdeal_Di@1 Vinm Vinp gnd net@23 Ideal_Differencer_1
XIdeal_Sa@0 Clock net@23 net@1 vdd Ideal_Sample_Hold
XIdeal_Sw@0 gnd net@1 vdd Vout Ideal_Switch
XIdeal_Sw@1 net@1 gnd Vout gnd Ideal_Switch
.ENDS Ideal_clocked_comparator

.global gnd vdd

*** TOP LEVEL CELL: Fig29_23_V2{sch}
Rres@0 Vout net@0 10000
Rres@1 net@2 gnd 1000
Rres@2 Vout net@8 10000
Rres@3 net@10 net@2 1000
Rres@4 Vout net@14 10000
Rres@5 net@16 net@10 1000
Rres@6 Vout net@20 10000
Rres@7 net@22 net@16 1000
Rres@8 Vout net@26 10000
Rres@9 net@28 net@22 1000
Rres@10 Vout net@32 10000
Rres@11 net@34 net@28 1000
Rres@12 Vout net@38 10000
Rres@13 net@40 net@34 1000
Rres@14 vdd net@129 1000
Rres@15 Vout gnd 10000
Rres@16 net@129 net@40 1000
Rres@17 net@129 net@40 1000
Rres@18 net@2 gnd 1000
XIdeal_cl@0 Vclock net@2 Vin net@0 vdd Ideal_clocked_comparator
XIdeal_cl@1 Vclock net@10 Vin net@8 vdd Ideal_clocked_comparator
XIdeal_cl@2 Vclock net@16 Vin net@14 vdd Ideal_clocked_comparator
XIdeal_cl@3 Vclock net@22 Vin net@20 vdd Ideal_clocked_comparator
XIdeal_cl@4 Vclock net@28 Vin net@26 vdd Ideal_clocked_comparator
XIdeal_cl@5 Vclock net@34 Vin net@32 vdd Ideal_clocked_comparator
XIdeal_cl@6 Vclock net@40 Vin net@38 vdd Ideal_clocked_comparator

* Spice Code nodes in cell cell 'Fig29_23_V2{sch}'
VDD VDD 0 DC 5
Vtrip Vtrip 0 DC 2.5
VGND GND 0 DC 0
Vin Vin 0 DC 0 PULSE(0 5 0 5u)
Vclock Vclock 0 DC 0 PULSE(0 5 5n 100p 100p 4.9n 10n)
.options post
.options plotwinsize=0
.tran 10p 5u 10p .1n uic
.END
