** Profile: "Fig9_30_PMOS-dc"  [ C:\Users\jbaker\Desktop\Chap9_PSpice\Fig9_30_PMOS\Fig9_30_pmos-pspicefiles\Fig9_30_pmos\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig9_30_pmos-pspicefiles/Fig9_30_pmos.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VSG 0 1 1m 
.TEMP 0 50 100
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig9_30_PMOS.net" 


.END
