** Profile: "Fig9_33_PMOS-dc"  [ C:\Users\jbaker\Desktop\Chap9_PSpice\Fig9_33_PMOS\Fig9_33_pmos-pspicefiles\Fig9_33_pmos\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig9_33_pmos-pspicefiles/Fig9_33_pmos.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VSG 0 500m 1m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig9_33_PMOS.net" 


.END
