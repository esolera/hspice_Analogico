*** Figure 29.3 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vout

*** CELL: Ideal_Switch{sch}
.SUBCKT Ideal_Switch contrlm contrlp in out

* Spice Code nodes in cell cell 'Ideal_Switch{sch}'
Sswitch  in out  contrlp contrlm  switmod
.model switmod sw
.ENDS Ideal_Switch

.global gnd vdd

*** TOP LEVEL CELL: Fig29_3{sch}
Rres@0 net@6 gnd 625
Rres@1 net@5 net@6 625
Rres@2 net@4 net@5 625
Rres@3 net@3 net@4 625
Rres@4 net@52 net@3 625
Rres@6 net@0 net@52 625
Rres@7 net@87 net@0 625
Rres@8 vdd net@87 625
XIdeal_Sw@0 Vtrip D0 net@6 A Ideal_Switch
XIdeal_Sw@1 Vtrip D0i net@5 net@15 Ideal_Switch
XIdeal_Sw@2 Vtrip D0 net@4 net@15 Ideal_Switch
XIdeal_Sw@3 Vtrip D0i net@3 net@23 Ideal_Switch
XIdeal_Sw@4 Vtrip D0 net@52 net@23 Ideal_Switch
XIdeal_Sw@5 Vtrip D0i net@0 net@31 Ideal_Switch
XIdeal_Sw@7 Vtrip D0i gnd A Ideal_Switch
XIdeal_Sw@8 Vtrip D0 net@87 net@31 Ideal_Switch
XIdeal_Sw@9 Vtrip D1 net@31 B Ideal_Switch
XIdeal_Sw@12 Vtrip D1i net@23 B Ideal_Switch
XIdeal_Sw@13 Vtrip D1 net@15 net@59 Ideal_Switch
XIdeal_Sw@14 Vtrip D1i A net@59 Ideal_Switch
XIdeal_Sw@15 Vtrip D2 B Vout Ideal_Switch
XIdeal_Sw@16 Vtrip D2i net@59 Vout Ideal_Switch

* Spice Code nodes in cell cell 'Fig29_3{sch}'
VDD VDD 0 DC 5
Vtrip Vtrip 0 DC 2.5
VGND GND 0 DC 0
VD0 D0 0 DC 0 PULSE(0 5 5n 100p 100p 4.9n 10n)
VD0i D0i 0 DC 0 PULSE(5 0  5n 100p 100p 4.9n 10n)
VD1 D1 0 DC 0 PULSE(0 5 10n 100p 100p 9.9n 20n)
VD1i D1i 0 DC 0 PULSE(5 0 10n 100p 100p 9.9n 20n)
VD2 D2 0 DC 0 PULSE(0 5 20n 100p 100p 19.9n 40n)
VD2i D2i 0 DC 0 PULSE(5 0 20n 100p 100p 19.9n 40n)
.options post
.options plotwinsize=0
.tran 10p 40n 10p .1n uic
.END
