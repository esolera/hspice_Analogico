*** Figure 1.11 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#print all

.op

Vin	Vin	0	DC	1
R1	Vin	Vout	1k
R2	Vout	0	2k

.end