*** Figure 24.24 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#set units=degrees
*#plot vout vin xlimit 400n 700n ylimit .4 1

.option scale=50n ITL1=300 vntol=1u abstol=1u reltol=1u
.tran 1n 700n UIC

VDD 	VDD	0	DC	1	

Vin	Vin	0	DC	0	PULSE 500m  900m 500n 0 0 50n 1u

Cc	Vout	Vd4t	240f
Cl	Vout	0	1000f

M1	vd1	vout	vss	0	N_50n L=2 W=50
M2	vout1	vin	vss	0	N_50n L=2 W=50
M6B	Vdb1	Vbias4	0	0	N_50n L=2 W=100
M6T	vss	Vbias3	vdb1	0	N_50n L=2 W=100
M3T	vd3t	vd1	VDD	VDD	P_50n L=1 W=100
M3B	vd1	vd1	vd3t	VDD	P_50n L=1 W=100
M4T	vd4t	vd1	VDD	VDD	P_50n L=1 W=100
M4B	vout1	vd1	vd4t	VDD	P_50n L=1 W=100


M7T	vd7t	Vout1	VDD	VDD	P_50n L=1 W=100
M7B	Vout	Vout1	vd7t	VDD	P_50n L=1 W=100

M8T	Vout	vbias3	vd8b	0	N_50n L=2 W=50
M8B	vd8b	vbias4	0	0	N_50n L=2 W=50


Xbias	VDD Vbias1 Vbias2 Vbias3 Vbias4 Vhigh Vlow Vncas Vpcas bias


.subckt bias VDD Vbias1 Vbias2 Vbias3 Vbias4 Vhigh Vlow Vncas Vpcas

MP1	Vbias3	Vbiasp	VDD	VDD	P_50n L=2 W=100
MP2	Vbias4	Vbiasp 	VDD	VDD	P_50n L=2 W=100
MP3	vp1	vp2	VDD	VDD	P_50n L=2 W=100
MP4	vp2	Vbias2	vp1	VDD	P_50n L=2 W=100
MP5	Vpcas	Vpcas	vp2	VDD	P_50n L=2 W=100
MP6	Vbias2	Vbias2	VDD	VDD	P_50n L=10 W=20
MP7	Vhigh	Vbias1	VDD	VDD	P_50n L=2 W=100
MP8	Vbias1	Vbias2	Vhigh	VDD	P_50n L=2 W=100
MP9	vp3	Vbias1	VDD	VDD	P_50n L=2 W=100
MP10	Vncas	Vbias2	vp3	VDD	P_50n L=2 W=100

MN1	Vbias3	Vbias3	0	0	N_50n L=10 W=10
MN2	Vbias4	Vbias3	Vlow	0	N_50n L=2 W=50
MN3	Vlow	Vbias4	0	0	N_50n L=2 W=50
MN4	Vpcas	Vbias3	vn1	0	N_50n L=2 W=50
MN5	vn1	Vbias4	0	0	N_50n L=2 W=50
MN6	Vbias2	Vbias3	vn2	0	N_50n L=2 W=50
MN7	vn2	Vbias4	0	0	N_50n L=2 W=50
MN8	Vbias1	Vbias3	vn3	0	N_50n L=2 W=50
MN9	vn3	Vbias4	0	0	N_50n L=2 W=50
MN10	Vncas	Vncas	vn4	0	N_50n L=2 W=50
MN11	vn4	Vbias3	vn5	0	N_50n L=2 W=50
MN12	vn5	vn4	0	0	N_50n L=2 W=50

MBM1	Vbiasn	Vbiasn	0	0	N_50n L=2 W=50
MBM2	Vreg	Vreg	Vr	0	N_50n L=2 W=200
MBM3	Vbiasn	Vbiasp	VDD	VDD	P_50n L=2 W=100
MBM4	Vreg	Vbiasp	VDD	VDD	P_50n L=2 W=100

Rbias	Vr	0	5.5k

*amplifier 
MA1	Vamp	Vreg	0	0	N_50n L=2 W=50
MA2	Vbiasp	Vbiasn	0	0	N_50n L=2 W=50
MA3	Vamp	Vamp	VDD	VDD	P_50n L=2 W=100
MA4	Vbiasp	Vamp	VDD	VDD	P_50n L=2 W=100

MCP	VDD	Vbiasp	VDD	VDD	P_50n L=100 W=100

*start-up stuff
MSU1	Vsur	Vbiasn	0	0	N_50n L=2   W=50
MSU2	Vsur	Vsur	VDD	VDD	P_50n L=20  W=10
MSU3	Vbiasp	Vsur	Vbiasn	0	N_50n L=1   W=10

.ends

.include cmosedu_models.txt 

.end
   

