*** Example 8.12 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot onoise_spectrum 
*#print all

.noise	V(Vout,0)	Vs 	dec  	100 	1 	100G 

Vs	Vs	0	dc	1.7	ac	1
Rs	Vs	Vout	1k
D1	Vout	0 	Diode

.model Diode D TT=10n Rs=0
.print noise all
.end