*** Figure 30.15 CMOS: Circuit Design, Layout, and Simulation ***

.tran 1n 3000n 10n 1n UIC

*#destroy all
*#run
*#plot Vout 

CL Vout 0 10p
VDD VDD 0 DC 1
VREFP VREFP 0 DC 1
VREFM VREFM 0 DC 0.0

VB9 B9 0 DC 0 pulse 1 0 0 200p 200p 1000n 2000n
VB8 B8 0 DC 0 
VB7 B7 0 DC 0 
VB6 B6 0 DC 1 
VB5 B5 0 DC 0 
VB4 B4 0 DC 0 
VB3 B3 0 DC 0 
VB2 B2 0 DC 0 
VB1 B1 0 DC 0 
VB0 B0 0 DC 0 

*Generate Logic switching point, or trip, voltage
R1 VDD trip 100MEG
R2 trip 0   100MEG

*Make resistive ladder
X9 trip B9 in9 Vout Vrefp Vrefm R2R
X8 trip B8 in8 in9 Vrefp Vrefm R2R
X7 trip B7 in7 in8 Vrefp Vrefm R2R
X6 trip B6 in6 in7 Vrefp Vrefm R2R
X5 trip B5 in5 in6 Vrefp Vrefm R2R
X4 trip B4 in4 in5 Vrefp Vrefm R2R
X3 trip B3 in3 in4 Vrefp Vrefm R2R
X2 trip B2 in2 in3 Vrefp Vrefm R2R
X1 trip B1 in1 in2 Vrefp Vrefm R2R
X0 trip B0 in0 in1 Vrefp Vrefm R2R
RT in0 0 10k

.subckt R2R trip BX in out Vrefp Vrefm
SH 	Vrefp	2R	BX	trip 	Switmod
SL	Vrefm	2R	trip	BX	Switmod
R2R	2R	out	20k
R1R	out	in	10k	
.model switmod SW
.ends

.end
