*** Figure 29.3_sine CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vout vin

VDD VDD 0 5
R1 VDD N001 625
R2 N001 N003 625
R3 N003 N005 625
R4 N005 N007 625
R5 N007 N008 625
R6 N008 N011 625
R7 N011 N013 625
R8 N013 0 625
XX1 N002 N001 D0 VDD switch_1
XX5 N002 N003 D0i VDD switch_1
XX6 N006 N005 D0 VDD switch_1
XX7 N006 N007 D0i VDD switch_1
XX8 N009 N008 D0 VDD switch_1
XX9 N009 N011 D0i VDD switch_1
XX10 N014 N013 D0 VDD switch_1
XX11 N014 0 D0i VDD switch_1
XX12 N004 N002 D1 VDD switch_1
XX13 N004 N006 D1i VDD switch_1
XX14 Vout N004 D2 VDD switch_1
XX15 N012 N009 D1 VDD switch_1
XX16 N012 N014 D1i VDD switch_1
XX17 Vout N012 D2i VDD switch_1
XX2 D2 D2i VDD inverter
XX3 D1 D1i VDD inverter
XX4 D0 D0i VDD inverter
Vclock1 N010 0 PULSE(0 5 5n 100p 100p 4.9n 10n)
Vin1 Vin 0 SINE(2.5 2 2MEG)
XX18 D2 D1 D0 Vin VDD 0 N010 VDD ideal_3_bit_adc

* block symbol definitions
.subckt switch_1 P1 P2 clk VDD
S1 P2 P1 clk Vtrip switmod
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
.model switmod SW
.ends switch_1

.subckt inverter In Out VDD
S3 Out VDD N001 In switmod
S4 0 Out In N001 switmod
E1 N001 0 VDD 0 0.5
.model switmod SW
.ends inverter

.subckt ideal_3_bit_adc B2 B1 B0 Vin Vrefp Vrefm Clock VDD
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
B1 VCM 0 V=(V(VREFP)-V(VREFM))/2
BPIP PIPIN 0 V=V(OUTSH)-V(VREFM)+((V(VREFP)-V(VREFM))/16)
XU7 VDD Vtrip VCM PIPIN B2 N001 adcbit
XU8 VDD Vtrip VCM N001 B1 N002 adcbit
XU9 VDD Vtrip VCM N002 B0 NC_01 adcbit
XU10 Vin OUTSH clock VDD sample_and_hold
.ends ideal_3_bit_adc

.subckt adcbit VDD Vtrip VCM Vin Bitout Vout
S3 Bitout VDD Vin VCM switmod
S4 0 Bitout VCM Vin switmod
S5 Vout Vinh Bitout Vtrip switmod
S6 Vinl Vout Vtrip Bitout switmod
E1 Vinh 0 Vin VCM 2
E2 Vinl 0 Vin 0 2
.model switmod SW
.ends adcbit

.subckt sample_and_hold Vin Outsh Clock VDD
S1 Vins Vinb Vtrip Clock switmod
C1 Vins 0 1e-10
S2 N001 Vins clock Vtrip switmod
C2 N001 0 1e-16
R1 Vtrip 0 100MEG
R2 VDD Vtrip 100MEG
Ebufout Outsh 0 N001 0 1
Ebufin Vinb 0 Vin 0 1
.model switmod SW
.ends sample_and_hold

.tran 0 2000n 0 .1n uic
.options plotwinsize=0

.end
