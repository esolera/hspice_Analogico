*** Figure 9.29 (PMOS) CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#set temp=0
*#run
*#set temp=50
*#run
*#set temp=100
*#run
*#plot -dc1.vsd#branch -dc2.vsd#branch -dc3.vsd#branch 

.option scale=1u
.DC 	VSG	0.8	1.8	1m

VSD 	0	VSD	DC	2
VSG	0	VSG	DC	0

M1	VSD	VSG	0	0	P_1u L=2 W=30
                                                                     
.include cmosedu_models.txt 

.end
      
