** Profile: "_Fig5_8_MSD-_Fig5_8_MSD"  [ C:\Users\Christian\Desktop\MSD\Ch5_MSD_PSpice\_Fig5_8_MSD\_Fig5_8_MSD-pspicefiles\_Fig5_8_MSD\_Fig5_8_MSD.sim ] 

** Creating circuit file "_Fig5_8_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 .01n 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig5_8_MSD.net" 


.END
