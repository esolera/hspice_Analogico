** Profile: "Fig10_12_PMOS_short-tran"  [ C:\Users\jbaker\Desktop\Chap10_PSpice\Fig10_12_PMOS_short\Fig10_12_pmos_short-pspicefiles\Fig10_12_pmos_short\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig10_12_pmos_short-pspicefiles/Fig10_12_pmos_short.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 800p 0 SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig10_12_PMOS_short.net" 


.END
