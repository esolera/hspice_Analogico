** Profile: "Fig10_12_NMOS_long-tran"  [ C:\Users\jbaker\Desktop\Chap10_PSpice\Fig10_12_NMOS_long\Fig10_12_nmos_long-pspicefiles\Fig10_12_nmos_long\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig10_12_nmos_long-pspicefiles/Fig10_12_nmos_long.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 600p 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig10_12_NMOS_long.net" 


.END
