** Profile: "Fig6_19_PMOS_ID_VSD-dc"  [ C:\USERS\STUDENT\DESKTOP\CHAP6_PSPICE\Fig6_19_PMOS_ID_VSD\Fig6_19_PMOS_ID_VSD-PSpiceFiles\Fig6_19_PMOS_ID_VSD\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../fig6_19_pmos_id_vsd-pspicefiles/fig6_19_pmos_id_vsd.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VSD 0 1 0.01 
+ LIN V_VSG 0 1 250m 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig6_19_PMOS_ID_VSD.net" 


.END
