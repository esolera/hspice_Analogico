*** Figure 28.10 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vout

*** CELL: Ideal_Switch{sch}
.SUBCKT Ideal_Switch contrlm contrlp in out

* Spice Code nodes in cell cell 'Ideal_Switch{sch}'
Sswitch  in out  contrlp contrlm  switmod
.model switmod sw
.ENDS Ideal_Switch

*** CELL: Ideal_DACbit{sch}
.SUBCKT Ideal_DACbit Bitin Bitout Vone Vtrip
** GLOBAL gnd
Xideal_sw@0 Bitin Vtrip Bitout gnd Ideal_Switch
Xideal_sw@1 Vtrip Bitin Vone Bitout Ideal_Switch
.ENDS Ideal_DACbit

*** CELL: Ideal_3Bit_DAC{sch}
.SUBCKT Ideal_3Bit_DAC B0 B1 B2 VREFM VREFP Vout vdd
** GLOBAL gnd
Rres@0 vdd Vtrip 100000k
Rres@1 Vtrip gnd 100000k
Rres@2 VREFP VREFM 100000k
XIdeal_DA@3 B2 B2L Vone Vtrip Ideal_DACbit
XIdeal_DA@6 B1 B1L Vone Vtrip Ideal_DACbit
XIdeal_DA@9 B0 B0L Vone Vtrip Ideal_DACbit

* Spice Code nodes in cell cell 'Ideal_3Bit_DAC{sch}'
Vone Vone 0 DC 1
B1 Vout 0 V=((v(vrefp)-v(vrefm))/8)*(v(B2L)*4+v(B1L)*2+v(B0L))+v(vrefm)
.ENDS Ideal_3Bit_DAC

.global gnd vdd

*** TOP LEVEL CELL: Fig28_10{sch}
XIdeal_3B@0 B0 B1 B2 gnd vdd Vout vdd Ideal_3Bit_DAC

* Spice Code nodes in cell cell 'Fig28_10{sch}'
VDD VDD 0 DC 1
VGND GND 0 DC 0
VB0 B0 0 DC 0 PULSE(0 1 5n 100p 100p 4.9n 10n)
VB1 B1 0 DC 0 PULSE(0 1 10n 100p 100p 9.9n 20n)
VB2 B2 0 DC 0 PULSE(0 1 20n 100p 100p 19.9n 40n)
.tran 10p 40n 10p .1n uic
.options post
.options plotwinsize=0
.END
