*** Figure 29.10 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot voutp voutm

*** CELL: Ideal_Switch{sch}
.SUBCKT Ideal_Switch contrlm contrlp in out

* Spice Code nodes in cell cell 'Ideal_Switch{sch}'
Sswitch  in out  contrlp contrlm  switmod
.model switmod sw
.ENDS Ideal_Switch

.global gnd vdd

*** TOP LEVEL CELL: Fig29_10{sch}
Rres@0 vdd Voutm 100000
Rres@1 vdd Voutp 100000
IDCCurren@6 net@668 gnd DC 40uA
IDCCurren@7 net@679 gnd DC 20uA
IDCCurren@8 net@718 gnd DC 10uA
XIdeal_Sw@16 Vtrip D2 Voutm net@668 Ideal_Switch
XIdeal_Sw@17 Vtrip D2i Voutp net@668 Ideal_Switch
XIdeal_Sw@18 Vtrip D1 Voutm net@679 Ideal_Switch
XIdeal_Sw@19 Vtrip D1i Voutp net@679 Ideal_Switch
XIdeal_Sw@20 Vtrip D0 Voutm net@718 Ideal_Switch
XIdeal_Sw@21 Vtrip D0i Voutp net@718 Ideal_Switch

* Spice Code nodes in cell cell 'Fig29_10{sch}'
VDD VDD 0 DC 5
Vtrip Vtrip 0 DC 2.5
VGND GND 0 DC 0
VD0 D0 0 DC 0 PULSE(0 5 5n 100p 100p 4.9n 10n)
VD0i D0i 0 DC 0 PULSE(5 0  5n 100p 100p 4.9n 10n)
VD1 D1 0 DC 0 PULSE(0 5 10n 100p 100p 9.9n 20n)
VD1i D1i 0 DC 0 PULSE(5 0 10n 100p 100p 9.9n 20n)
VD2 D2 0 DC 0 PULSE(0 5 20n 100p 100p 19.9n 40n)
VD2i D2i 0 DC 0 PULSE(5 0 20n 100p 100p 19.9n 40n)
.options post
.options plotwinsize=0
.tran 10p 40n 10p .1n uic
.END
