*** Figure 9.34 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#let ID=mag(VDS#branch)
*#let IG=mag(VGS#branch)
*#plot 20*log(ID/IG)


.option scale=50n
.AC	DEC 100	10MEG 10G

VDS 	VDS	0	DC	1
VGS	VGS	0	DC	350m	AC	1

M1	VDS	VGS	0	0	N_50n L=2 W=50

.include cmosedu_models.txt

.end
   
