** Profile: "_Fig3_46_MSD-_Fig3_46_MSD"  [ C:\Users\jbaker\Desktop\Ch3_MSD_PSpice\_fig3_46_msd-pspicefiles\_fig3_46_msd\_fig3_46_msd.sim ] 

** Creating circuit file "_Fig3_46_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1k 100meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig3_46_MSD.net" 


.END
