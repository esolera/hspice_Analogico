*** Example 8.5 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot onoise_spectrum
*#print all

.noise	 v(2,0)	vin dec  100 1 1k 
R1	 1 2 10k 
R2	 2 0 1k 
Vin	 1 0	dc 0 ac 1
.print noise all
.end