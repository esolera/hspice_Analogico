*** Figure 9.33 (PMOS) CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#let ID=-VSD#branch
*#let gm=deriv(ID)
*#plot gm


.option scale=50n
.DC 	VSG	0	500m	1m

VSD 	0	VSD	DC	100m
VSG	0	VSG	DC	0

M1	VSD	VSG	0	0	P_50n L=2 W=100

.include cmosedu_models.txt

.end
   
