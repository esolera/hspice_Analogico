*** Figure 3.7 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vin vout

.tran 1p 250p 

O1	Vin	0	Vout	0	TRC
Rload	Vout	0	1G
Vin	vin	0	DC	0	pulse 0 1 50p 0

.model TRC 	ltra	R=0.1 	C=32e-18 len=5000

.end
