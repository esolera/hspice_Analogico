*** Figure 26.4 CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot v:xbias:Vmeas1#branch
*#plot vbiasn vbiasp

.option scale=50n
.dc VDD 0 1.2 1m

VDD 	VDD	0	DC	1 pulse 0 1 100u

Xbias	vbiasn	vbiasp	VDD	bias

.subckt bias vbiasn vbiasp VDD

Vmeas1	Vmeas1	0	DC	0

M1	Vbiasn	Vbiasn	0	0	N_50n L=1 W=10
M2	Vreg	Vreg	Vr	0	N_50n L=1 W=40
M3	Vbiasn	Vbiasp	VDD	VDD	P_50n L=1 W=20
M4	Vreg	Vbiasp	VDD	VDD	P_50n L=1 W=20

Rbias	Vr	vmeas1	4k

*amplifier 
MA1	Vamp	Vreg	0	0	N_50n L=2 W=10
MA2	Vbiasp	Vbiasn	0	0	N_50n L=2 W=10
MA3	Vamp	Vamp	VDD	VDD	P_50n L=2 W=20
MA4	Vbiasp	Vamp	VDD	VDD	P_50n L=2 W=20

*start-up stuff
MSU1	Vsur	Vbiasn	0	0	N_50n L=1   W=10
MSU2	Vsur	Vsur	VDD	VDD	P_50n L=20  W=10
MSU3	Vbiasp	Vsur	Vbiasn	0	N_50n L=1   W=10

.ends

* 50nm BSIM4 models
*
* Don't forget the .options scale=50nm if using an Lmin of 1 
* 1<Ldrawn<200   10<Wdrawn<10000 Vdd=1V
* Change to level=54 when using HSPICE

.include cmosedu_models.txt

.end
   

