** Profile: "SCHEMATIC1-_Fig3_37_MSD"  [ C:\Users\HomePC\Documents\Spring 2013\PSpice_CMOSedu\MSD\Ch3_MSD_Pspice\_Fig3_37_MSD\_fig3_37_msd-pspicefiles\schematic1\_fig3_37_msd.sim ] 

** Creating circuit file "_Fig3_37_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 10k 100meg
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
