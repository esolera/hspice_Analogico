** Profile: "Fig6_12-DC Sweep"  [ C:\Users\student\Desktop\Chap6_PSpice\Fig6_12\Fig6_12-PSpiceFiles\Fig6_12\DC Sweep.sim ] 

** Creating circuit file "DC Sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../fig6_12-pspicefiles/fig6_12.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN VDS 0 5 0.01 
+ LIN VGS 0 5 1 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig6_12.net" 


.END
