** Profile: "Fig10_19_PMOS-tran"  [ C:\Users\jbaker\Desktop\Chap10_PSpice\Fig10_19_PMOS\Fig10_19_pmos-pspicefiles\Fig10_19_pmos\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig10_19_pmos-pspicefiles/Fig10_19_pmos.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2.5n 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig10_19_PMOS.net" 


.END
