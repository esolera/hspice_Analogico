*** Figure 26.1_nmos CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vgn 

.option scale=50n 
.dc	Idn	0	250u 	10n

VDD	VDD	0	DC	1

Idn	VDD	vgn	DC	0
**Idp	vgp	0	DC	0

Mn	vgn	vgn	0	0	N_50n L=1 W=10
**Mp	vgp	vgp	VDD	VDD	P_50n L=1 W=20

* 50nm BSIM4 models
*
* Don't forget the .options scale=50nm if using an Lmin of 1 
* 1<Ldrawn<200   10<Wdrawn<10000 Vdd=1V
* Change to level=54 when using HSPICE

.include cmosedu_models.txt

.end
   

