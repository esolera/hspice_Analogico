** Profile: "SCHEMATIC1-_Fig3_51_MSD"  [ C:\Users\HomePC\Desktop\MSD\Ch3_MSD_Pspice\_Fig3_51_MSD\_fig3_51_msd-pspicefiles\schematic1\_fig3_51_msd.sim ] 

** Creating circuit file "_Fig3_51_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 80u 0 .01u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
