** Profile: "Fig10_12_NMOS_short-tran"  [ C:\Users\jbaker\Desktop\Chap10_PSpice\Fig10_12_NMOS_short\Fig10_12_nmos_short-pspicefiles\Fig10_12_nmos_short\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig10_12_nmos_short-pspicefiles/Fig10_12_nmos_short.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1n 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig10_12_NMOS_short.net" 


.END
