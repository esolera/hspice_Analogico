** Profile: "NOISE_NMOS_50n-noise"  [ C:\Users\jbaker\Desktop\Chap9_PSpice\NOISE_NMOS_50n\Noise_nmos_50n-pspicefiles\Noise_nmos_50n\Noise.sim ] 

** Creating circuit file "noise.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Noise_nmos_50n-pspicefiles/Noise_nmos_50n.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 1000MEG
.NOISE V([VD],[0]) V_VGS 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\NOISE_NMOS_50n.net" 


.END
