** Profile: "Fig6_13_PMOS-dc"  [ C:\Users\jbaker\Desktop\PSpice_CMOSedu\Chap6_PSpice\Fig6_13_PMOS\Fig6_13_pmos-pspicefiles\Fig6_13_pmos\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../Fig6_13_pmos-pspicefiles/Fig6_13_pmos.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_VSG 0 2 1m 
+ LIN V_VBS 0 5 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Fig6_13_PMOS.net" 


.END
