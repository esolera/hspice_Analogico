** Profile: "_Fig2_18_MSD-_Fig2_18_MSD"  [ C:\Users\jbaker\Desktop\Ch2_MSD\_Fig2_18_MSD-pspicefiles\_Fig2_18_MSD\_Fig2_18_MSD.sim ] 

** Creating circuit file "_Fig2_18_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2us 0 .001us SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig2_18_MSD.net" 


.END
