** Profile: "_Fig3_49_MSD-_Fig3_49_MSD"  [ C:\Users\jbaker\Desktop\Ch3_MSD_PSpice\_Fig3_49_MSD-pspicefiles\_Fig3_49_MSD\_Fig3_49_MSD.sim ] 

** Creating circuit file "_Fig3_49_MSD.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10u 8u SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\_Fig3_49_MSD.net" 


.END
