*** Figure 28.5b CMOS: Circuit Design, Layout, and Simulation ***

*#destroy all
*#run
*#plot vin vout

*** CELL: Ideal_Switch{sch}
.SUBCKT Ideal_Switch contrlm contrlp in out

* Spice Code nodes in cell cell 'Ideal_Switch{sch}'
Sswitch  in out  contrlp contrlm  switmod
.model switmod sw
.ENDS Ideal_Switch

*** CELL: Ideal_Opamp{sch}
.SUBCKT Ideal_Opamp Vm Vo Vp
** GLOBAL gnd
Rres@0 Vp Vm 1410.065meg
Rres@1 Vo gnd 1

* Spice Code nodes in cell cell 'Ideal_Opamp{sch}'
G1 Vo 0  Vp  Vm 100MEG
.ENDS Ideal_Opamp

*** CELL: Ideal_Track&Hold{sch}
.SUBCKT Ideal_Track_Hold Vclk Vin Voutsh vdd
** GLOBAL gnd
Ccap@0 gnd Vins 0.1n
Rres@0 vdd Vtrip 100000k
Rres@1 Vtrip gnd 100000k
XIdeal_sw@0 Vclk Vtrip Vinb Vins Ideal_Switch
Xideal_op@0 Voutsh Voutsh Vins Ideal_Opamp
Xideal_op@1 Vinb Vinb Vin Ideal_Opamp
.ENDS Ideal_Track_Hold

.global gnd

*** TOP LEVEL CELL: Fig28_5b{sch}
XIdeal_Sa@0 Vclk Vin Vout vdd Ideal_Track_Hold

* Spice Code nodes in cell cell 'Fig28_5b{sch}'
VDD VDD 0 DC 1
VGND GND 0 DC 0
Vin Vin 0 DC 0 SINE(0.5 0.5 4MEG)
Vclk Vclk 0 DC 0 PULSE(0 1 0 0 0 4.9n 10n)
.tran 10p 500n 10p .1n
.options post
.options plotwinsize=0
.END
